module efm_lut_decoder
(
  input   [13:0] i_efm_symb,
  output  [7:0]  o_data,
  
  output         o_s0_sync,
  output         o_s1_sync
);

reg [7:0] r_data;
assign o_data = r_data;
assign o_s0_sync = i_efm_symb == 14'b00100000000001;
assign o_s1_sync = i_efm_symb == 14'b00000000010010;

always@(*) begin
  case(i_efm_symb)
    14'b01001000100000: r_data <= 8'd0  ;
    14'b10000100000000: r_data <= 8'd1  ;
    14'b10010000100000: r_data <= 8'd2  ;
    14'b10001000100000: r_data <= 8'd3  ;
    14'b01000100000000: r_data <= 8'd4  ;
    14'b00000100010000: r_data <= 8'd5  ;
    14'b00010000100000: r_data <= 8'd6  ;
    14'b00100100000000: r_data <= 8'd7  ;
    14'b01001001000000: r_data <= 8'd8  ;
    14'b10000001000000: r_data <= 8'd9  ;
    14'b10010001000000: r_data <= 8'd10 ;
    14'b10001001000000: r_data <= 8'd11 ;
    14'b01000001000000: r_data <= 8'd12 ;
    14'b00000001000000: r_data <= 8'd13 ;
    14'b00010001000000: r_data <= 8'd14 ;
    14'b00100001000000: r_data <= 8'd15 ;
    14'b10000000100000: r_data <= 8'd16 ;
    14'b10000010000000: r_data <= 8'd17 ;
    14'b10010010000000: r_data <= 8'd18 ;
    14'b00100000100000: r_data <= 8'd19 ;
    14'b01000010000000: r_data <= 8'd20 ;
    14'b00000010000000: r_data <= 8'd21 ;
    14'b00010010000000: r_data <= 8'd22 ;
    14'b00100010000000: r_data <= 8'd23 ;
    14'b01001000010000: r_data <= 8'd24 ;
    14'b10000000010000: r_data <= 8'd25 ;
    14'b10010000010000: r_data <= 8'd26 ;
    14'b10001000010000: r_data <= 8'd27 ;
    14'b01000000010000: r_data <= 8'd28 ;
    14'b00001000010000: r_data <= 8'd29 ;
    14'b00010000010000: r_data <= 8'd30 ;
    14'b00100000010000: r_data <= 8'd31 ;
    14'b00000000100000: r_data <= 8'd32 ;
    14'b10000100001000: r_data <= 8'd33 ;
    14'b00001000100000: r_data <= 8'd34 ;
    14'b00100100100000: r_data <= 8'd35 ;
    14'b01000100001000: r_data <= 8'd36 ;
    14'b00000100001000: r_data <= 8'd37 ;
    14'b01000000100000: r_data <= 8'd38 ;
    14'b00100100001000: r_data <= 8'd39 ;
    14'b01001001001000: r_data <= 8'd40 ;
    14'b10000001001000: r_data <= 8'd41 ;
    14'b10010001001000: r_data <= 8'd42 ;
    14'b10001001001000: r_data <= 8'd43 ;
    14'b01000001001000: r_data <= 8'd44 ;
    14'b00000001001000: r_data <= 8'd45 ;
    14'b00010001001000: r_data <= 8'd46 ;
    14'b00100001001000: r_data <= 8'd47 ;
    14'b00000100000000: r_data <= 8'd48 ;
    14'b10000010001000: r_data <= 8'd49 ;
    14'b10010010001000: r_data <= 8'd50 ;
    14'b10000100010000: r_data <= 8'd51 ;
    14'b01000010001000: r_data <= 8'd52 ;
    14'b00000010001000: r_data <= 8'd53 ;
    14'b00010010001000: r_data <= 8'd54 ;
    14'b00100010001000: r_data <= 8'd55 ;
    14'b01001000001000: r_data <= 8'd56 ;
    14'b10000000001000: r_data <= 8'd57 ;
    14'b10010000001000: r_data <= 8'd58 ;
    14'b10001000001000: r_data <= 8'd59 ;
    14'b01000000001000: r_data <= 8'd60 ;
    14'b00001000001000: r_data <= 8'd61 ;
    14'b00010000001000: r_data <= 8'd62 ;
    14'b00100000001000: r_data <= 8'd63 ;
    14'b01001000100100: r_data <= 8'd64 ;
    14'b10000100100100: r_data <= 8'd65 ;
    14'b10010000100100: r_data <= 8'd66 ;
    14'b10001000100100: r_data <= 8'd67 ;
    14'b01000100100100: r_data <= 8'd68 ;
    14'b00000000100100: r_data <= 8'd69 ;
    14'b00010000100100: r_data <= 8'd70 ;
    14'b00100100100100: r_data <= 8'd71 ;
    14'b01001001000100: r_data <= 8'd72 ;
    14'b10000001000100: r_data <= 8'd73 ;
    14'b10010001000100: r_data <= 8'd74 ;
    14'b10001001000100: r_data <= 8'd75 ;
    14'b01000001000100: r_data <= 8'd76 ;
    14'b00000001000100: r_data <= 8'd77 ;
    14'b00010001000100: r_data <= 8'd78 ;
    14'b00100001000100: r_data <= 8'd79 ;
    14'b10000000100100: r_data <= 8'd80 ;
    14'b10000010000100: r_data <= 8'd81 ;
    14'b10010010000100: r_data <= 8'd82 ;
    14'b00100000100100: r_data <= 8'd83 ;
    14'b01000010000100: r_data <= 8'd84 ;
    14'b00000010000100: r_data <= 8'd85 ;
    14'b00010010000100: r_data <= 8'd86 ;
    14'b00100010000100: r_data <= 8'd87 ;
    14'b01001000000100: r_data <= 8'd88 ;
    14'b10000000000100: r_data <= 8'd89 ;
    14'b10010000000100: r_data <= 8'd90 ;
    14'b10001000000100: r_data <= 8'd91 ;
    14'b01000000000100: r_data <= 8'd92 ;
    14'b00001000000100: r_data <= 8'd93 ;
    14'b00010000000100: r_data <= 8'd94 ;
    14'b00100000000100: r_data <= 8'd95 ;
    14'b01001000100010: r_data <= 8'd96 ;
    14'b10000100100010: r_data <= 8'd97 ;
    14'b10010000100010: r_data <= 8'd98 ;
    14'b10001000100010: r_data <= 8'd99 ;
    14'b01000100100010: r_data <= 8'd100;
    14'b00000000100010: r_data <= 8'd101;
    14'b01000000100100: r_data <= 8'd102;
    14'b00100100100010: r_data <= 8'd103;
    14'b01001001000010: r_data <= 8'd104;
    14'b10000001000010: r_data <= 8'd105;
    14'b10010001000010: r_data <= 8'd106;
    14'b10001001000010: r_data <= 8'd107;
    14'b01000001000010: r_data <= 8'd108;
    14'b00000001000010: r_data <= 8'd109;
    14'b00010001000010: r_data <= 8'd110;
    14'b00100001000010: r_data <= 8'd111;
    14'b10000000100010: r_data <= 8'd112;
    14'b10000010000010: r_data <= 8'd113;
    14'b10010010000010: r_data <= 8'd114;
    14'b00100000100010: r_data <= 8'd115;
    14'b01000010000010: r_data <= 8'd116;
    14'b00000010000010: r_data <= 8'd117;
    14'b00010010000010: r_data <= 8'd118;
    14'b00100010000010: r_data <= 8'd119;
    14'b01001000000010: r_data <= 8'd120;
    14'b00001001001000: r_data <= 8'd121;
    14'b10010000000010: r_data <= 8'd122;
    14'b10001000000010: r_data <= 8'd123;
    14'b01000000000010: r_data <= 8'd124;
    14'b00001000000010: r_data <= 8'd125;
    14'b00010000000010: r_data <= 8'd126;
    14'b00100000000010: r_data <= 8'd127;
    14'b01001000100001: r_data <= 8'd128;
    14'b10000100100001: r_data <= 8'd129;
    14'b10010000100001: r_data <= 8'd130;
    14'b10001000100001: r_data <= 8'd131;
    14'b01000100100001: r_data <= 8'd132;
    14'b00000000100001: r_data <= 8'd133;
    14'b00010000100001: r_data <= 8'd134;
    14'b00100100100001: r_data <= 8'd135;
    14'b01001001000001: r_data <= 8'd136;
    14'b10000001000001: r_data <= 8'd137;
    14'b10010001000001: r_data <= 8'd138;
    14'b10001001000001: r_data <= 8'd139;
    14'b01000001000001: r_data <= 8'd140;
    14'b00000001000001: r_data <= 8'd141;
    14'b00010001000001: r_data <= 8'd142;
    14'b00100001000001: r_data <= 8'd143;
    14'b10000000100001: r_data <= 8'd144;
    14'b10000010000001: r_data <= 8'd145;
    14'b10010010000001: r_data <= 8'd146;
    14'b00100000100001: r_data <= 8'd147;
    14'b01000010000001: r_data <= 8'd148;
    14'b00000010000001: r_data <= 8'd149;
    14'b00010010000001: r_data <= 8'd150;
    14'b00100010000001: r_data <= 8'd151;
    14'b01001000000001: r_data <= 8'd152;
    14'b10000010010000: r_data <= 8'd153;
    14'b10010000000001: r_data <= 8'd154;
    14'b10001000000001: r_data <= 8'd155;
    14'b01000010010000: r_data <= 8'd156;
    14'b00001000000001: r_data <= 8'd157;
    14'b00010000000001: r_data <= 8'd158;
    14'b00100010010000: r_data <= 8'd159;
    14'b00001000100001: r_data <= 8'd160;
    14'b10000100001001: r_data <= 8'd161;
    14'b01000100010000: r_data <= 8'd162;
    14'b00000100100001: r_data <= 8'd163;
    14'b01000100001001: r_data <= 8'd164;
    14'b00000100001001: r_data <= 8'd165;
    14'b01000000100001: r_data <= 8'd166;
    14'b00100100001001: r_data <= 8'd167;
    14'b01001001001001: r_data <= 8'd168;
    14'b10000001001001: r_data <= 8'd169;
    14'b10010001001001: r_data <= 8'd170;
    14'b10001001001001: r_data <= 8'd171;
    14'b01000001001001: r_data <= 8'd172;
    14'b00000001001001: r_data <= 8'd173;
    14'b00010001001001: r_data <= 8'd174;
    14'b00100001001001: r_data <= 8'd175;
    14'b00000100100000: r_data <= 8'd176;
    14'b10000010001001: r_data <= 8'd177;
    14'b10010010001001: r_data <= 8'd178;
    14'b00100100010000: r_data <= 8'd179;
    14'b01000010001001: r_data <= 8'd180;
    14'b00000010001001: r_data <= 8'd181;
    14'b00010010001001: r_data <= 8'd182;
    14'b00100010001001: r_data <= 8'd183;
    14'b01001000001001: r_data <= 8'd184;
    14'b10000000001001: r_data <= 8'd185;
    14'b10010000001001: r_data <= 8'd186;
    14'b10001000001001: r_data <= 8'd187;
    14'b01000000001001: r_data <= 8'd188;
    14'b00001000001001: r_data <= 8'd189;
    14'b00010000001001: r_data <= 8'd190;
    14'b00100000001001: r_data <= 8'd191;
    14'b01000100100000: r_data <= 8'd192;
    14'b10000100010001: r_data <= 8'd193;
    14'b10010010010000: r_data <= 8'd194;
    14'b00001000100100: r_data <= 8'd195;
    14'b01000100010001: r_data <= 8'd196;
    14'b00000100010001: r_data <= 8'd197;
    14'b00010010010000: r_data <= 8'd198;
    14'b00100100010001: r_data <= 8'd199;
    14'b00001001000001: r_data <= 8'd200;
    14'b10000100000001: r_data <= 8'd201;
    14'b00001001000100: r_data <= 8'd202;
    14'b00001001000000: r_data <= 8'd203;
    14'b01000100000001: r_data <= 8'd204;
    14'b00000100000001: r_data <= 8'd205;
    14'b00000010010000: r_data <= 8'd206;
    14'b00100100000001: r_data <= 8'd207;
    14'b00000100100100: r_data <= 8'd208;
    14'b10000010010001: r_data <= 8'd209;
    14'b10010010010001: r_data <= 8'd210;
    14'b10000100100000: r_data <= 8'd211;
    14'b01000010010001: r_data <= 8'd212;
    14'b00000010010001: r_data <= 8'd213;
    14'b00010010010001: r_data <= 8'd214;
    14'b00100010010001: r_data <= 8'd215;
    14'b01001000010001: r_data <= 8'd216;
    14'b10000000010001: r_data <= 8'd217;
    14'b10010000010001: r_data <= 8'd218;
    14'b10001000010001: r_data <= 8'd219;
    14'b01000000010001: r_data <= 8'd220;
    14'b00001000010001: r_data <= 8'd221;
    14'b00010000010001: r_data <= 8'd222;
    14'b00100000010001: r_data <= 8'd223;
    14'b01000100000010: r_data <= 8'd224;
    14'b00000100000010: r_data <= 8'd225;
    14'b10000100010010: r_data <= 8'd226;
    14'b00100100000010: r_data <= 8'd227;
    14'b01000100010010: r_data <= 8'd228;
    14'b00000100010010: r_data <= 8'd229;
    14'b01000000100010: r_data <= 8'd230;
    14'b00100100010010: r_data <= 8'd231;
    14'b10000100000010: r_data <= 8'd232;
    14'b10000100000100: r_data <= 8'd233;
    14'b00001001001001: r_data <= 8'd234;
    14'b00001001000010: r_data <= 8'd235;
    14'b01000100000100: r_data <= 8'd236;
    14'b00000100000100: r_data <= 8'd237;
    14'b00010000100010: r_data <= 8'd238;
    14'b00100100000100: r_data <= 8'd239;
    14'b00000100100010: r_data <= 8'd240;
    14'b10000010010010: r_data <= 8'd241;
    14'b10010010010010: r_data <= 8'd242;
    14'b00001000100010: r_data <= 8'd243;
    14'b01000010010010: r_data <= 8'd244;
    14'b00000010010010: r_data <= 8'd245;
    14'b00010010010010: r_data <= 8'd246;
    14'b00100010010010: r_data <= 8'd247;
    14'b01001000010010: r_data <= 8'd248;
    14'b10000000010010: r_data <= 8'd249;
    14'b10010000010010: r_data <= 8'd250;
    14'b10001000010010: r_data <= 8'd251;
    14'b01000000010010: r_data <= 8'd252;
    14'b00001000010010: r_data <= 8'd253;
    14'b00010000010010: r_data <= 8'd254;
    14'b00100000010010: r_data <= 8'd255;
	default: r_data <= 8'd0;
  endcase
end
endmodule
