// GF(256) multiplier + accumulator
// Vladislav Knyazkov, October 2023

module gf256_mac(
    input [7:0] a,
    input [7:0] b,
    input [7:0] c,

    output [7:0] s
);

endmodule
